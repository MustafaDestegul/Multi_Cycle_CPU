module Producer7(out7,out0);
output reg [2:0] out7;
output reg [2:0] out0;




always 
begin 
	out7<=3'd7;
	out0<=3'd2;
end



endmodule
