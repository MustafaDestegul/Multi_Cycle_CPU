module RandomNumberGenerator(out);
output reg [7:0] out;




always 
begin 
	out<=8'b00001111;
end



endmodule
