module Producer0(out);
output reg [7:0] out;




always 
begin 
	out<=8'd0;
end



endmodule
