module producer4(out);
output reg [7:0] out;




always 
begin 
	out<=8'd4;
end



endmodule
